class hello;

  function new();
    // Nothing to do here
  endfunction

  function void print_hello();
    $display("Hello, World");
  endfunction

endclass
